module control_unit(
output reg	Gra, Grb, Grc, RIn, ROut, BAOut, CONin,
				HiIn, LoIn, ZIn, PCIn, MDRIn, MARIn, YIn, OPortIn, IRIn,
				HiOut, LoOut, ZHiOut, ZLoOut, PCOut, MDROut, IPortOut, COut,
				Read, Write, Clear, Run,
output reg[4:0] ALUCode,
input[31:0] IR,
input			Clock, Reset, Stop, CON_FF

);


endmodule