module RAM (
	input wire r, w, //active high
	input wire [8:0] addr,
	input wire [31:0] din,
	output reg [31:0] dout,
	input wire START
);


reg [31:0] mem [0:511];

always @(*) begin
		dout <= 32'b0;
	if(r == 1) begin
		dout <= mem[addr];
	end else if(w == 1) begin
		mem[addr] <= din;
	end
	if(START == 1) begin
	mem['h54] = 'h97;//for ld instructions
 mem['hDB] = 'h46;

//3.1.1 ld R4, 0x54;
 mem[32'd311] = 32'b_00000_0100_0000_00000000000_01010100;

//3.1.2 ld R6, 0x63(R2);
 mem[32'd312] = 32'b_00000_0110_0010_00000000000_01100011;

//3.1.3 ldi R4, 0x54;
 mem[32'd313] = 32'b_00001_0100_0000_00000000000_01010100;

//3.1.4 ldi R6, 0x63(R2);
 mem[32'd314] = 32'b_00001_0110_0010_00000000000_01100011;



 mem['h34] = 'h25;//for st instructions
 mem['hEA] = 'h19;

//3.2.1 st 0x34, R3;
 mem[32'd321] = 32'b00010_0011_0000_00000000000_00110100;

//3.2.2 st 0x34(R3), R3;
 mem[32'd322] = 32'b00010_0011_0011_00000000000_00110100;

 
 
//3.3.1 addi R5, R6, -7;
 mem[32'd331] = 32'b01100_0101_0110_11111111111_11111001;
//3.3.2 andi R5, R6, 0x95;
 mem[32'd332] = 32'b01100_0101_0110_00000000000_10010101;

//3.3.3 ori R5, R6, 0x95;
 mem[32'd333] = 32'b01110_0101_0110_00000000000_10010101;



//3.4.1 brzr R1, 27;
 mem[32'd341] = 32'b10011_0001_0000_00000000000_00011011;

//3.4.2 brnz R1, 27;
 mem[32'd342] = 32'b10011_0001_0001_00000000000_00011011;

//3.4.3 brpl R1, 27;
 mem[32'd343] = 32'b10011_0001_0010_00000000000_00011011;

//3.4.4 brmi R1, 27;
 mem[32'd344] = 32'b10011_0001_0011_00000000000_00011011;



//3.5.1 jr R8;
 mem[32'd351] = 32'b10101_1000_0000_00000000000_00000000;

//3.5.2 jal R5;
 mem[32'd352] = 32'b10100_0101_1000_00000000000_00000000;



//3.6.1 mfhi R3
 mem[32'd361] = 32'b11001_0011_0000_00000000000_00000000;
//3.6.2 mflo R2
 mem[32'd362] = 32'b11000_0010_0000_00000000000_00000000;



//3.7.1 out R6
 mem[32'd371] = 32'b10110_0110_0000_00000000000_00000000;
//3.7.2 in R3
 mem[32'd372] = 32'b10111_0011_0000_00000000000_00000000;
 end
end

endmodule